-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: ula_mux.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.0.0 Build 614 04/24/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY ula_mux IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END ula_mux;


ARCHITECTURE SYN OF ula_mux IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (20 DOWNTO 0, 31 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
	sub_wire21    <= data0x(31 DOWNTO 0);
	sub_wire20    <= data1x(31 DOWNTO 0);
	sub_wire19    <= data2x(31 DOWNTO 0);
	sub_wire18    <= data3x(31 DOWNTO 0);
	sub_wire17    <= data4x(31 DOWNTO 0);
	sub_wire16    <= data5x(31 DOWNTO 0);
	sub_wire15    <= data6x(31 DOWNTO 0);
	sub_wire14    <= data7x(31 DOWNTO 0);
	sub_wire13    <= data8x(31 DOWNTO 0);
	sub_wire12    <= data9x(31 DOWNTO 0);
	sub_wire11    <= data10x(31 DOWNTO 0);
	sub_wire10    <= data11x(31 DOWNTO 0);
	sub_wire9    <= data12x(31 DOWNTO 0);
	sub_wire8    <= data13x(31 DOWNTO 0);
	sub_wire7    <= data14x(31 DOWNTO 0);
	sub_wire6    <= data15x(31 DOWNTO 0);
	sub_wire5    <= data16x(31 DOWNTO 0);
	sub_wire4    <= data17x(31 DOWNTO 0);
	sub_wire3    <= data18x(31 DOWNTO 0);
	sub_wire2    <= data19x(31 DOWNTO 0);
	sub_wire0    <= data20x(31 DOWNTO 0);
	sub_wire1(20, 0)    <= sub_wire0(0);
	sub_wire1(20, 1)    <= sub_wire0(1);
	sub_wire1(20, 2)    <= sub_wire0(2);
	sub_wire1(20, 3)    <= sub_wire0(3);
	sub_wire1(20, 4)    <= sub_wire0(4);
	sub_wire1(20, 5)    <= sub_wire0(5);
	sub_wire1(20, 6)    <= sub_wire0(6);
	sub_wire1(20, 7)    <= sub_wire0(7);
	sub_wire1(20, 8)    <= sub_wire0(8);
	sub_wire1(20, 9)    <= sub_wire0(9);
	sub_wire1(20, 10)    <= sub_wire0(10);
	sub_wire1(20, 11)    <= sub_wire0(11);
	sub_wire1(20, 12)    <= sub_wire0(12);
	sub_wire1(20, 13)    <= sub_wire0(13);
	sub_wire1(20, 14)    <= sub_wire0(14);
	sub_wire1(20, 15)    <= sub_wire0(15);
	sub_wire1(20, 16)    <= sub_wire0(16);
	sub_wire1(20, 17)    <= sub_wire0(17);
	sub_wire1(20, 18)    <= sub_wire0(18);
	sub_wire1(20, 19)    <= sub_wire0(19);
	sub_wire1(20, 20)    <= sub_wire0(20);
	sub_wire1(20, 21)    <= sub_wire0(21);
	sub_wire1(20, 22)    <= sub_wire0(22);
	sub_wire1(20, 23)    <= sub_wire0(23);
	sub_wire1(20, 24)    <= sub_wire0(24);
	sub_wire1(20, 25)    <= sub_wire0(25);
	sub_wire1(20, 26)    <= sub_wire0(26);
	sub_wire1(20, 27)    <= sub_wire0(27);
	sub_wire1(20, 28)    <= sub_wire0(28);
	sub_wire1(20, 29)    <= sub_wire0(29);
	sub_wire1(20, 30)    <= sub_wire0(30);
	sub_wire1(20, 31)    <= sub_wire0(31);
	sub_wire1(19, 0)    <= sub_wire2(0);
	sub_wire1(19, 1)    <= sub_wire2(1);
	sub_wire1(19, 2)    <= sub_wire2(2);
	sub_wire1(19, 3)    <= sub_wire2(3);
	sub_wire1(19, 4)    <= sub_wire2(4);
	sub_wire1(19, 5)    <= sub_wire2(5);
	sub_wire1(19, 6)    <= sub_wire2(6);
	sub_wire1(19, 7)    <= sub_wire2(7);
	sub_wire1(19, 8)    <= sub_wire2(8);
	sub_wire1(19, 9)    <= sub_wire2(9);
	sub_wire1(19, 10)    <= sub_wire2(10);
	sub_wire1(19, 11)    <= sub_wire2(11);
	sub_wire1(19, 12)    <= sub_wire2(12);
	sub_wire1(19, 13)    <= sub_wire2(13);
	sub_wire1(19, 14)    <= sub_wire2(14);
	sub_wire1(19, 15)    <= sub_wire2(15);
	sub_wire1(19, 16)    <= sub_wire2(16);
	sub_wire1(19, 17)    <= sub_wire2(17);
	sub_wire1(19, 18)    <= sub_wire2(18);
	sub_wire1(19, 19)    <= sub_wire2(19);
	sub_wire1(19, 20)    <= sub_wire2(20);
	sub_wire1(19, 21)    <= sub_wire2(21);
	sub_wire1(19, 22)    <= sub_wire2(22);
	sub_wire1(19, 23)    <= sub_wire2(23);
	sub_wire1(19, 24)    <= sub_wire2(24);
	sub_wire1(19, 25)    <= sub_wire2(25);
	sub_wire1(19, 26)    <= sub_wire2(26);
	sub_wire1(19, 27)    <= sub_wire2(27);
	sub_wire1(19, 28)    <= sub_wire2(28);
	sub_wire1(19, 29)    <= sub_wire2(29);
	sub_wire1(19, 30)    <= sub_wire2(30);
	sub_wire1(19, 31)    <= sub_wire2(31);
	sub_wire1(18, 0)    <= sub_wire3(0);
	sub_wire1(18, 1)    <= sub_wire3(1);
	sub_wire1(18, 2)    <= sub_wire3(2);
	sub_wire1(18, 3)    <= sub_wire3(3);
	sub_wire1(18, 4)    <= sub_wire3(4);
	sub_wire1(18, 5)    <= sub_wire3(5);
	sub_wire1(18, 6)    <= sub_wire3(6);
	sub_wire1(18, 7)    <= sub_wire3(7);
	sub_wire1(18, 8)    <= sub_wire3(8);
	sub_wire1(18, 9)    <= sub_wire3(9);
	sub_wire1(18, 10)    <= sub_wire3(10);
	sub_wire1(18, 11)    <= sub_wire3(11);
	sub_wire1(18, 12)    <= sub_wire3(12);
	sub_wire1(18, 13)    <= sub_wire3(13);
	sub_wire1(18, 14)    <= sub_wire3(14);
	sub_wire1(18, 15)    <= sub_wire3(15);
	sub_wire1(18, 16)    <= sub_wire3(16);
	sub_wire1(18, 17)    <= sub_wire3(17);
	sub_wire1(18, 18)    <= sub_wire3(18);
	sub_wire1(18, 19)    <= sub_wire3(19);
	sub_wire1(18, 20)    <= sub_wire3(20);
	sub_wire1(18, 21)    <= sub_wire3(21);
	sub_wire1(18, 22)    <= sub_wire3(22);
	sub_wire1(18, 23)    <= sub_wire3(23);
	sub_wire1(18, 24)    <= sub_wire3(24);
	sub_wire1(18, 25)    <= sub_wire3(25);
	sub_wire1(18, 26)    <= sub_wire3(26);
	sub_wire1(18, 27)    <= sub_wire3(27);
	sub_wire1(18, 28)    <= sub_wire3(28);
	sub_wire1(18, 29)    <= sub_wire3(29);
	sub_wire1(18, 30)    <= sub_wire3(30);
	sub_wire1(18, 31)    <= sub_wire3(31);
	sub_wire1(17, 0)    <= sub_wire4(0);
	sub_wire1(17, 1)    <= sub_wire4(1);
	sub_wire1(17, 2)    <= sub_wire4(2);
	sub_wire1(17, 3)    <= sub_wire4(3);
	sub_wire1(17, 4)    <= sub_wire4(4);
	sub_wire1(17, 5)    <= sub_wire4(5);
	sub_wire1(17, 6)    <= sub_wire4(6);
	sub_wire1(17, 7)    <= sub_wire4(7);
	sub_wire1(17, 8)    <= sub_wire4(8);
	sub_wire1(17, 9)    <= sub_wire4(9);
	sub_wire1(17, 10)    <= sub_wire4(10);
	sub_wire1(17, 11)    <= sub_wire4(11);
	sub_wire1(17, 12)    <= sub_wire4(12);
	sub_wire1(17, 13)    <= sub_wire4(13);
	sub_wire1(17, 14)    <= sub_wire4(14);
	sub_wire1(17, 15)    <= sub_wire4(15);
	sub_wire1(17, 16)    <= sub_wire4(16);
	sub_wire1(17, 17)    <= sub_wire4(17);
	sub_wire1(17, 18)    <= sub_wire4(18);
	sub_wire1(17, 19)    <= sub_wire4(19);
	sub_wire1(17, 20)    <= sub_wire4(20);
	sub_wire1(17, 21)    <= sub_wire4(21);
	sub_wire1(17, 22)    <= sub_wire4(22);
	sub_wire1(17, 23)    <= sub_wire4(23);
	sub_wire1(17, 24)    <= sub_wire4(24);
	sub_wire1(17, 25)    <= sub_wire4(25);
	sub_wire1(17, 26)    <= sub_wire4(26);
	sub_wire1(17, 27)    <= sub_wire4(27);
	sub_wire1(17, 28)    <= sub_wire4(28);
	sub_wire1(17, 29)    <= sub_wire4(29);
	sub_wire1(17, 30)    <= sub_wire4(30);
	sub_wire1(17, 31)    <= sub_wire4(31);
	sub_wire1(16, 0)    <= sub_wire5(0);
	sub_wire1(16, 1)    <= sub_wire5(1);
	sub_wire1(16, 2)    <= sub_wire5(2);
	sub_wire1(16, 3)    <= sub_wire5(3);
	sub_wire1(16, 4)    <= sub_wire5(4);
	sub_wire1(16, 5)    <= sub_wire5(5);
	sub_wire1(16, 6)    <= sub_wire5(6);
	sub_wire1(16, 7)    <= sub_wire5(7);
	sub_wire1(16, 8)    <= sub_wire5(8);
	sub_wire1(16, 9)    <= sub_wire5(9);
	sub_wire1(16, 10)    <= sub_wire5(10);
	sub_wire1(16, 11)    <= sub_wire5(11);
	sub_wire1(16, 12)    <= sub_wire5(12);
	sub_wire1(16, 13)    <= sub_wire5(13);
	sub_wire1(16, 14)    <= sub_wire5(14);
	sub_wire1(16, 15)    <= sub_wire5(15);
	sub_wire1(16, 16)    <= sub_wire5(16);
	sub_wire1(16, 17)    <= sub_wire5(17);
	sub_wire1(16, 18)    <= sub_wire5(18);
	sub_wire1(16, 19)    <= sub_wire5(19);
	sub_wire1(16, 20)    <= sub_wire5(20);
	sub_wire1(16, 21)    <= sub_wire5(21);
	sub_wire1(16, 22)    <= sub_wire5(22);
	sub_wire1(16, 23)    <= sub_wire5(23);
	sub_wire1(16, 24)    <= sub_wire5(24);
	sub_wire1(16, 25)    <= sub_wire5(25);
	sub_wire1(16, 26)    <= sub_wire5(26);
	sub_wire1(16, 27)    <= sub_wire5(27);
	sub_wire1(16, 28)    <= sub_wire5(28);
	sub_wire1(16, 29)    <= sub_wire5(29);
	sub_wire1(16, 30)    <= sub_wire5(30);
	sub_wire1(16, 31)    <= sub_wire5(31);
	sub_wire1(15, 0)    <= sub_wire6(0);
	sub_wire1(15, 1)    <= sub_wire6(1);
	sub_wire1(15, 2)    <= sub_wire6(2);
	sub_wire1(15, 3)    <= sub_wire6(3);
	sub_wire1(15, 4)    <= sub_wire6(4);
	sub_wire1(15, 5)    <= sub_wire6(5);
	sub_wire1(15, 6)    <= sub_wire6(6);
	sub_wire1(15, 7)    <= sub_wire6(7);
	sub_wire1(15, 8)    <= sub_wire6(8);
	sub_wire1(15, 9)    <= sub_wire6(9);
	sub_wire1(15, 10)    <= sub_wire6(10);
	sub_wire1(15, 11)    <= sub_wire6(11);
	sub_wire1(15, 12)    <= sub_wire6(12);
	sub_wire1(15, 13)    <= sub_wire6(13);
	sub_wire1(15, 14)    <= sub_wire6(14);
	sub_wire1(15, 15)    <= sub_wire6(15);
	sub_wire1(15, 16)    <= sub_wire6(16);
	sub_wire1(15, 17)    <= sub_wire6(17);
	sub_wire1(15, 18)    <= sub_wire6(18);
	sub_wire1(15, 19)    <= sub_wire6(19);
	sub_wire1(15, 20)    <= sub_wire6(20);
	sub_wire1(15, 21)    <= sub_wire6(21);
	sub_wire1(15, 22)    <= sub_wire6(22);
	sub_wire1(15, 23)    <= sub_wire6(23);
	sub_wire1(15, 24)    <= sub_wire6(24);
	sub_wire1(15, 25)    <= sub_wire6(25);
	sub_wire1(15, 26)    <= sub_wire6(26);
	sub_wire1(15, 27)    <= sub_wire6(27);
	sub_wire1(15, 28)    <= sub_wire6(28);
	sub_wire1(15, 29)    <= sub_wire6(29);
	sub_wire1(15, 30)    <= sub_wire6(30);
	sub_wire1(15, 31)    <= sub_wire6(31);
	sub_wire1(14, 0)    <= sub_wire7(0);
	sub_wire1(14, 1)    <= sub_wire7(1);
	sub_wire1(14, 2)    <= sub_wire7(2);
	sub_wire1(14, 3)    <= sub_wire7(3);
	sub_wire1(14, 4)    <= sub_wire7(4);
	sub_wire1(14, 5)    <= sub_wire7(5);
	sub_wire1(14, 6)    <= sub_wire7(6);
	sub_wire1(14, 7)    <= sub_wire7(7);
	sub_wire1(14, 8)    <= sub_wire7(8);
	sub_wire1(14, 9)    <= sub_wire7(9);
	sub_wire1(14, 10)    <= sub_wire7(10);
	sub_wire1(14, 11)    <= sub_wire7(11);
	sub_wire1(14, 12)    <= sub_wire7(12);
	sub_wire1(14, 13)    <= sub_wire7(13);
	sub_wire1(14, 14)    <= sub_wire7(14);
	sub_wire1(14, 15)    <= sub_wire7(15);
	sub_wire1(14, 16)    <= sub_wire7(16);
	sub_wire1(14, 17)    <= sub_wire7(17);
	sub_wire1(14, 18)    <= sub_wire7(18);
	sub_wire1(14, 19)    <= sub_wire7(19);
	sub_wire1(14, 20)    <= sub_wire7(20);
	sub_wire1(14, 21)    <= sub_wire7(21);
	sub_wire1(14, 22)    <= sub_wire7(22);
	sub_wire1(14, 23)    <= sub_wire7(23);
	sub_wire1(14, 24)    <= sub_wire7(24);
	sub_wire1(14, 25)    <= sub_wire7(25);
	sub_wire1(14, 26)    <= sub_wire7(26);
	sub_wire1(14, 27)    <= sub_wire7(27);
	sub_wire1(14, 28)    <= sub_wire7(28);
	sub_wire1(14, 29)    <= sub_wire7(29);
	sub_wire1(14, 30)    <= sub_wire7(30);
	sub_wire1(14, 31)    <= sub_wire7(31);
	sub_wire1(13, 0)    <= sub_wire8(0);
	sub_wire1(13, 1)    <= sub_wire8(1);
	sub_wire1(13, 2)    <= sub_wire8(2);
	sub_wire1(13, 3)    <= sub_wire8(3);
	sub_wire1(13, 4)    <= sub_wire8(4);
	sub_wire1(13, 5)    <= sub_wire8(5);
	sub_wire1(13, 6)    <= sub_wire8(6);
	sub_wire1(13, 7)    <= sub_wire8(7);
	sub_wire1(13, 8)    <= sub_wire8(8);
	sub_wire1(13, 9)    <= sub_wire8(9);
	sub_wire1(13, 10)    <= sub_wire8(10);
	sub_wire1(13, 11)    <= sub_wire8(11);
	sub_wire1(13, 12)    <= sub_wire8(12);
	sub_wire1(13, 13)    <= sub_wire8(13);
	sub_wire1(13, 14)    <= sub_wire8(14);
	sub_wire1(13, 15)    <= sub_wire8(15);
	sub_wire1(13, 16)    <= sub_wire8(16);
	sub_wire1(13, 17)    <= sub_wire8(17);
	sub_wire1(13, 18)    <= sub_wire8(18);
	sub_wire1(13, 19)    <= sub_wire8(19);
	sub_wire1(13, 20)    <= sub_wire8(20);
	sub_wire1(13, 21)    <= sub_wire8(21);
	sub_wire1(13, 22)    <= sub_wire8(22);
	sub_wire1(13, 23)    <= sub_wire8(23);
	sub_wire1(13, 24)    <= sub_wire8(24);
	sub_wire1(13, 25)    <= sub_wire8(25);
	sub_wire1(13, 26)    <= sub_wire8(26);
	sub_wire1(13, 27)    <= sub_wire8(27);
	sub_wire1(13, 28)    <= sub_wire8(28);
	sub_wire1(13, 29)    <= sub_wire8(29);
	sub_wire1(13, 30)    <= sub_wire8(30);
	sub_wire1(13, 31)    <= sub_wire8(31);
	sub_wire1(12, 0)    <= sub_wire9(0);
	sub_wire1(12, 1)    <= sub_wire9(1);
	sub_wire1(12, 2)    <= sub_wire9(2);
	sub_wire1(12, 3)    <= sub_wire9(3);
	sub_wire1(12, 4)    <= sub_wire9(4);
	sub_wire1(12, 5)    <= sub_wire9(5);
	sub_wire1(12, 6)    <= sub_wire9(6);
	sub_wire1(12, 7)    <= sub_wire9(7);
	sub_wire1(12, 8)    <= sub_wire9(8);
	sub_wire1(12, 9)    <= sub_wire9(9);
	sub_wire1(12, 10)    <= sub_wire9(10);
	sub_wire1(12, 11)    <= sub_wire9(11);
	sub_wire1(12, 12)    <= sub_wire9(12);
	sub_wire1(12, 13)    <= sub_wire9(13);
	sub_wire1(12, 14)    <= sub_wire9(14);
	sub_wire1(12, 15)    <= sub_wire9(15);
	sub_wire1(12, 16)    <= sub_wire9(16);
	sub_wire1(12, 17)    <= sub_wire9(17);
	sub_wire1(12, 18)    <= sub_wire9(18);
	sub_wire1(12, 19)    <= sub_wire9(19);
	sub_wire1(12, 20)    <= sub_wire9(20);
	sub_wire1(12, 21)    <= sub_wire9(21);
	sub_wire1(12, 22)    <= sub_wire9(22);
	sub_wire1(12, 23)    <= sub_wire9(23);
	sub_wire1(12, 24)    <= sub_wire9(24);
	sub_wire1(12, 25)    <= sub_wire9(25);
	sub_wire1(12, 26)    <= sub_wire9(26);
	sub_wire1(12, 27)    <= sub_wire9(27);
	sub_wire1(12, 28)    <= sub_wire9(28);
	sub_wire1(12, 29)    <= sub_wire9(29);
	sub_wire1(12, 30)    <= sub_wire9(30);
	sub_wire1(12, 31)    <= sub_wire9(31);
	sub_wire1(11, 0)    <= sub_wire10(0);
	sub_wire1(11, 1)    <= sub_wire10(1);
	sub_wire1(11, 2)    <= sub_wire10(2);
	sub_wire1(11, 3)    <= sub_wire10(3);
	sub_wire1(11, 4)    <= sub_wire10(4);
	sub_wire1(11, 5)    <= sub_wire10(5);
	sub_wire1(11, 6)    <= sub_wire10(6);
	sub_wire1(11, 7)    <= sub_wire10(7);
	sub_wire1(11, 8)    <= sub_wire10(8);
	sub_wire1(11, 9)    <= sub_wire10(9);
	sub_wire1(11, 10)    <= sub_wire10(10);
	sub_wire1(11, 11)    <= sub_wire10(11);
	sub_wire1(11, 12)    <= sub_wire10(12);
	sub_wire1(11, 13)    <= sub_wire10(13);
	sub_wire1(11, 14)    <= sub_wire10(14);
	sub_wire1(11, 15)    <= sub_wire10(15);
	sub_wire1(11, 16)    <= sub_wire10(16);
	sub_wire1(11, 17)    <= sub_wire10(17);
	sub_wire1(11, 18)    <= sub_wire10(18);
	sub_wire1(11, 19)    <= sub_wire10(19);
	sub_wire1(11, 20)    <= sub_wire10(20);
	sub_wire1(11, 21)    <= sub_wire10(21);
	sub_wire1(11, 22)    <= sub_wire10(22);
	sub_wire1(11, 23)    <= sub_wire10(23);
	sub_wire1(11, 24)    <= sub_wire10(24);
	sub_wire1(11, 25)    <= sub_wire10(25);
	sub_wire1(11, 26)    <= sub_wire10(26);
	sub_wire1(11, 27)    <= sub_wire10(27);
	sub_wire1(11, 28)    <= sub_wire10(28);
	sub_wire1(11, 29)    <= sub_wire10(29);
	sub_wire1(11, 30)    <= sub_wire10(30);
	sub_wire1(11, 31)    <= sub_wire10(31);
	sub_wire1(10, 0)    <= sub_wire11(0);
	sub_wire1(10, 1)    <= sub_wire11(1);
	sub_wire1(10, 2)    <= sub_wire11(2);
	sub_wire1(10, 3)    <= sub_wire11(3);
	sub_wire1(10, 4)    <= sub_wire11(4);
	sub_wire1(10, 5)    <= sub_wire11(5);
	sub_wire1(10, 6)    <= sub_wire11(6);
	sub_wire1(10, 7)    <= sub_wire11(7);
	sub_wire1(10, 8)    <= sub_wire11(8);
	sub_wire1(10, 9)    <= sub_wire11(9);
	sub_wire1(10, 10)    <= sub_wire11(10);
	sub_wire1(10, 11)    <= sub_wire11(11);
	sub_wire1(10, 12)    <= sub_wire11(12);
	sub_wire1(10, 13)    <= sub_wire11(13);
	sub_wire1(10, 14)    <= sub_wire11(14);
	sub_wire1(10, 15)    <= sub_wire11(15);
	sub_wire1(10, 16)    <= sub_wire11(16);
	sub_wire1(10, 17)    <= sub_wire11(17);
	sub_wire1(10, 18)    <= sub_wire11(18);
	sub_wire1(10, 19)    <= sub_wire11(19);
	sub_wire1(10, 20)    <= sub_wire11(20);
	sub_wire1(10, 21)    <= sub_wire11(21);
	sub_wire1(10, 22)    <= sub_wire11(22);
	sub_wire1(10, 23)    <= sub_wire11(23);
	sub_wire1(10, 24)    <= sub_wire11(24);
	sub_wire1(10, 25)    <= sub_wire11(25);
	sub_wire1(10, 26)    <= sub_wire11(26);
	sub_wire1(10, 27)    <= sub_wire11(27);
	sub_wire1(10, 28)    <= sub_wire11(28);
	sub_wire1(10, 29)    <= sub_wire11(29);
	sub_wire1(10, 30)    <= sub_wire11(30);
	sub_wire1(10, 31)    <= sub_wire11(31);
	sub_wire1(9, 0)    <= sub_wire12(0);
	sub_wire1(9, 1)    <= sub_wire12(1);
	sub_wire1(9, 2)    <= sub_wire12(2);
	sub_wire1(9, 3)    <= sub_wire12(3);
	sub_wire1(9, 4)    <= sub_wire12(4);
	sub_wire1(9, 5)    <= sub_wire12(5);
	sub_wire1(9, 6)    <= sub_wire12(6);
	sub_wire1(9, 7)    <= sub_wire12(7);
	sub_wire1(9, 8)    <= sub_wire12(8);
	sub_wire1(9, 9)    <= sub_wire12(9);
	sub_wire1(9, 10)    <= sub_wire12(10);
	sub_wire1(9, 11)    <= sub_wire12(11);
	sub_wire1(9, 12)    <= sub_wire12(12);
	sub_wire1(9, 13)    <= sub_wire12(13);
	sub_wire1(9, 14)    <= sub_wire12(14);
	sub_wire1(9, 15)    <= sub_wire12(15);
	sub_wire1(9, 16)    <= sub_wire12(16);
	sub_wire1(9, 17)    <= sub_wire12(17);
	sub_wire1(9, 18)    <= sub_wire12(18);
	sub_wire1(9, 19)    <= sub_wire12(19);
	sub_wire1(9, 20)    <= sub_wire12(20);
	sub_wire1(9, 21)    <= sub_wire12(21);
	sub_wire1(9, 22)    <= sub_wire12(22);
	sub_wire1(9, 23)    <= sub_wire12(23);
	sub_wire1(9, 24)    <= sub_wire12(24);
	sub_wire1(9, 25)    <= sub_wire12(25);
	sub_wire1(9, 26)    <= sub_wire12(26);
	sub_wire1(9, 27)    <= sub_wire12(27);
	sub_wire1(9, 28)    <= sub_wire12(28);
	sub_wire1(9, 29)    <= sub_wire12(29);
	sub_wire1(9, 30)    <= sub_wire12(30);
	sub_wire1(9, 31)    <= sub_wire12(31);
	sub_wire1(8, 0)    <= sub_wire13(0);
	sub_wire1(8, 1)    <= sub_wire13(1);
	sub_wire1(8, 2)    <= sub_wire13(2);
	sub_wire1(8, 3)    <= sub_wire13(3);
	sub_wire1(8, 4)    <= sub_wire13(4);
	sub_wire1(8, 5)    <= sub_wire13(5);
	sub_wire1(8, 6)    <= sub_wire13(6);
	sub_wire1(8, 7)    <= sub_wire13(7);
	sub_wire1(8, 8)    <= sub_wire13(8);
	sub_wire1(8, 9)    <= sub_wire13(9);
	sub_wire1(8, 10)    <= sub_wire13(10);
	sub_wire1(8, 11)    <= sub_wire13(11);
	sub_wire1(8, 12)    <= sub_wire13(12);
	sub_wire1(8, 13)    <= sub_wire13(13);
	sub_wire1(8, 14)    <= sub_wire13(14);
	sub_wire1(8, 15)    <= sub_wire13(15);
	sub_wire1(8, 16)    <= sub_wire13(16);
	sub_wire1(8, 17)    <= sub_wire13(17);
	sub_wire1(8, 18)    <= sub_wire13(18);
	sub_wire1(8, 19)    <= sub_wire13(19);
	sub_wire1(8, 20)    <= sub_wire13(20);
	sub_wire1(8, 21)    <= sub_wire13(21);
	sub_wire1(8, 22)    <= sub_wire13(22);
	sub_wire1(8, 23)    <= sub_wire13(23);
	sub_wire1(8, 24)    <= sub_wire13(24);
	sub_wire1(8, 25)    <= sub_wire13(25);
	sub_wire1(8, 26)    <= sub_wire13(26);
	sub_wire1(8, 27)    <= sub_wire13(27);
	sub_wire1(8, 28)    <= sub_wire13(28);
	sub_wire1(8, 29)    <= sub_wire13(29);
	sub_wire1(8, 30)    <= sub_wire13(30);
	sub_wire1(8, 31)    <= sub_wire13(31);
	sub_wire1(7, 0)    <= sub_wire14(0);
	sub_wire1(7, 1)    <= sub_wire14(1);
	sub_wire1(7, 2)    <= sub_wire14(2);
	sub_wire1(7, 3)    <= sub_wire14(3);
	sub_wire1(7, 4)    <= sub_wire14(4);
	sub_wire1(7, 5)    <= sub_wire14(5);
	sub_wire1(7, 6)    <= sub_wire14(6);
	sub_wire1(7, 7)    <= sub_wire14(7);
	sub_wire1(7, 8)    <= sub_wire14(8);
	sub_wire1(7, 9)    <= sub_wire14(9);
	sub_wire1(7, 10)    <= sub_wire14(10);
	sub_wire1(7, 11)    <= sub_wire14(11);
	sub_wire1(7, 12)    <= sub_wire14(12);
	sub_wire1(7, 13)    <= sub_wire14(13);
	sub_wire1(7, 14)    <= sub_wire14(14);
	sub_wire1(7, 15)    <= sub_wire14(15);
	sub_wire1(7, 16)    <= sub_wire14(16);
	sub_wire1(7, 17)    <= sub_wire14(17);
	sub_wire1(7, 18)    <= sub_wire14(18);
	sub_wire1(7, 19)    <= sub_wire14(19);
	sub_wire1(7, 20)    <= sub_wire14(20);
	sub_wire1(7, 21)    <= sub_wire14(21);
	sub_wire1(7, 22)    <= sub_wire14(22);
	sub_wire1(7, 23)    <= sub_wire14(23);
	sub_wire1(7, 24)    <= sub_wire14(24);
	sub_wire1(7, 25)    <= sub_wire14(25);
	sub_wire1(7, 26)    <= sub_wire14(26);
	sub_wire1(7, 27)    <= sub_wire14(27);
	sub_wire1(7, 28)    <= sub_wire14(28);
	sub_wire1(7, 29)    <= sub_wire14(29);
	sub_wire1(7, 30)    <= sub_wire14(30);
	sub_wire1(7, 31)    <= sub_wire14(31);
	sub_wire1(6, 0)    <= sub_wire15(0);
	sub_wire1(6, 1)    <= sub_wire15(1);
	sub_wire1(6, 2)    <= sub_wire15(2);
	sub_wire1(6, 3)    <= sub_wire15(3);
	sub_wire1(6, 4)    <= sub_wire15(4);
	sub_wire1(6, 5)    <= sub_wire15(5);
	sub_wire1(6, 6)    <= sub_wire15(6);
	sub_wire1(6, 7)    <= sub_wire15(7);
	sub_wire1(6, 8)    <= sub_wire15(8);
	sub_wire1(6, 9)    <= sub_wire15(9);
	sub_wire1(6, 10)    <= sub_wire15(10);
	sub_wire1(6, 11)    <= sub_wire15(11);
	sub_wire1(6, 12)    <= sub_wire15(12);
	sub_wire1(6, 13)    <= sub_wire15(13);
	sub_wire1(6, 14)    <= sub_wire15(14);
	sub_wire1(6, 15)    <= sub_wire15(15);
	sub_wire1(6, 16)    <= sub_wire15(16);
	sub_wire1(6, 17)    <= sub_wire15(17);
	sub_wire1(6, 18)    <= sub_wire15(18);
	sub_wire1(6, 19)    <= sub_wire15(19);
	sub_wire1(6, 20)    <= sub_wire15(20);
	sub_wire1(6, 21)    <= sub_wire15(21);
	sub_wire1(6, 22)    <= sub_wire15(22);
	sub_wire1(6, 23)    <= sub_wire15(23);
	sub_wire1(6, 24)    <= sub_wire15(24);
	sub_wire1(6, 25)    <= sub_wire15(25);
	sub_wire1(6, 26)    <= sub_wire15(26);
	sub_wire1(6, 27)    <= sub_wire15(27);
	sub_wire1(6, 28)    <= sub_wire15(28);
	sub_wire1(6, 29)    <= sub_wire15(29);
	sub_wire1(6, 30)    <= sub_wire15(30);
	sub_wire1(6, 31)    <= sub_wire15(31);
	sub_wire1(5, 0)    <= sub_wire16(0);
	sub_wire1(5, 1)    <= sub_wire16(1);
	sub_wire1(5, 2)    <= sub_wire16(2);
	sub_wire1(5, 3)    <= sub_wire16(3);
	sub_wire1(5, 4)    <= sub_wire16(4);
	sub_wire1(5, 5)    <= sub_wire16(5);
	sub_wire1(5, 6)    <= sub_wire16(6);
	sub_wire1(5, 7)    <= sub_wire16(7);
	sub_wire1(5, 8)    <= sub_wire16(8);
	sub_wire1(5, 9)    <= sub_wire16(9);
	sub_wire1(5, 10)    <= sub_wire16(10);
	sub_wire1(5, 11)    <= sub_wire16(11);
	sub_wire1(5, 12)    <= sub_wire16(12);
	sub_wire1(5, 13)    <= sub_wire16(13);
	sub_wire1(5, 14)    <= sub_wire16(14);
	sub_wire1(5, 15)    <= sub_wire16(15);
	sub_wire1(5, 16)    <= sub_wire16(16);
	sub_wire1(5, 17)    <= sub_wire16(17);
	sub_wire1(5, 18)    <= sub_wire16(18);
	sub_wire1(5, 19)    <= sub_wire16(19);
	sub_wire1(5, 20)    <= sub_wire16(20);
	sub_wire1(5, 21)    <= sub_wire16(21);
	sub_wire1(5, 22)    <= sub_wire16(22);
	sub_wire1(5, 23)    <= sub_wire16(23);
	sub_wire1(5, 24)    <= sub_wire16(24);
	sub_wire1(5, 25)    <= sub_wire16(25);
	sub_wire1(5, 26)    <= sub_wire16(26);
	sub_wire1(5, 27)    <= sub_wire16(27);
	sub_wire1(5, 28)    <= sub_wire16(28);
	sub_wire1(5, 29)    <= sub_wire16(29);
	sub_wire1(5, 30)    <= sub_wire16(30);
	sub_wire1(5, 31)    <= sub_wire16(31);
	sub_wire1(4, 0)    <= sub_wire17(0);
	sub_wire1(4, 1)    <= sub_wire17(1);
	sub_wire1(4, 2)    <= sub_wire17(2);
	sub_wire1(4, 3)    <= sub_wire17(3);
	sub_wire1(4, 4)    <= sub_wire17(4);
	sub_wire1(4, 5)    <= sub_wire17(5);
	sub_wire1(4, 6)    <= sub_wire17(6);
	sub_wire1(4, 7)    <= sub_wire17(7);
	sub_wire1(4, 8)    <= sub_wire17(8);
	sub_wire1(4, 9)    <= sub_wire17(9);
	sub_wire1(4, 10)    <= sub_wire17(10);
	sub_wire1(4, 11)    <= sub_wire17(11);
	sub_wire1(4, 12)    <= sub_wire17(12);
	sub_wire1(4, 13)    <= sub_wire17(13);
	sub_wire1(4, 14)    <= sub_wire17(14);
	sub_wire1(4, 15)    <= sub_wire17(15);
	sub_wire1(4, 16)    <= sub_wire17(16);
	sub_wire1(4, 17)    <= sub_wire17(17);
	sub_wire1(4, 18)    <= sub_wire17(18);
	sub_wire1(4, 19)    <= sub_wire17(19);
	sub_wire1(4, 20)    <= sub_wire17(20);
	sub_wire1(4, 21)    <= sub_wire17(21);
	sub_wire1(4, 22)    <= sub_wire17(22);
	sub_wire1(4, 23)    <= sub_wire17(23);
	sub_wire1(4, 24)    <= sub_wire17(24);
	sub_wire1(4, 25)    <= sub_wire17(25);
	sub_wire1(4, 26)    <= sub_wire17(26);
	sub_wire1(4, 27)    <= sub_wire17(27);
	sub_wire1(4, 28)    <= sub_wire17(28);
	sub_wire1(4, 29)    <= sub_wire17(29);
	sub_wire1(4, 30)    <= sub_wire17(30);
	sub_wire1(4, 31)    <= sub_wire17(31);
	sub_wire1(3, 0)    <= sub_wire18(0);
	sub_wire1(3, 1)    <= sub_wire18(1);
	sub_wire1(3, 2)    <= sub_wire18(2);
	sub_wire1(3, 3)    <= sub_wire18(3);
	sub_wire1(3, 4)    <= sub_wire18(4);
	sub_wire1(3, 5)    <= sub_wire18(5);
	sub_wire1(3, 6)    <= sub_wire18(6);
	sub_wire1(3, 7)    <= sub_wire18(7);
	sub_wire1(3, 8)    <= sub_wire18(8);
	sub_wire1(3, 9)    <= sub_wire18(9);
	sub_wire1(3, 10)    <= sub_wire18(10);
	sub_wire1(3, 11)    <= sub_wire18(11);
	sub_wire1(3, 12)    <= sub_wire18(12);
	sub_wire1(3, 13)    <= sub_wire18(13);
	sub_wire1(3, 14)    <= sub_wire18(14);
	sub_wire1(3, 15)    <= sub_wire18(15);
	sub_wire1(3, 16)    <= sub_wire18(16);
	sub_wire1(3, 17)    <= sub_wire18(17);
	sub_wire1(3, 18)    <= sub_wire18(18);
	sub_wire1(3, 19)    <= sub_wire18(19);
	sub_wire1(3, 20)    <= sub_wire18(20);
	sub_wire1(3, 21)    <= sub_wire18(21);
	sub_wire1(3, 22)    <= sub_wire18(22);
	sub_wire1(3, 23)    <= sub_wire18(23);
	sub_wire1(3, 24)    <= sub_wire18(24);
	sub_wire1(3, 25)    <= sub_wire18(25);
	sub_wire1(3, 26)    <= sub_wire18(26);
	sub_wire1(3, 27)    <= sub_wire18(27);
	sub_wire1(3, 28)    <= sub_wire18(28);
	sub_wire1(3, 29)    <= sub_wire18(29);
	sub_wire1(3, 30)    <= sub_wire18(30);
	sub_wire1(3, 31)    <= sub_wire18(31);
	sub_wire1(2, 0)    <= sub_wire19(0);
	sub_wire1(2, 1)    <= sub_wire19(1);
	sub_wire1(2, 2)    <= sub_wire19(2);
	sub_wire1(2, 3)    <= sub_wire19(3);
	sub_wire1(2, 4)    <= sub_wire19(4);
	sub_wire1(2, 5)    <= sub_wire19(5);
	sub_wire1(2, 6)    <= sub_wire19(6);
	sub_wire1(2, 7)    <= sub_wire19(7);
	sub_wire1(2, 8)    <= sub_wire19(8);
	sub_wire1(2, 9)    <= sub_wire19(9);
	sub_wire1(2, 10)    <= sub_wire19(10);
	sub_wire1(2, 11)    <= sub_wire19(11);
	sub_wire1(2, 12)    <= sub_wire19(12);
	sub_wire1(2, 13)    <= sub_wire19(13);
	sub_wire1(2, 14)    <= sub_wire19(14);
	sub_wire1(2, 15)    <= sub_wire19(15);
	sub_wire1(2, 16)    <= sub_wire19(16);
	sub_wire1(2, 17)    <= sub_wire19(17);
	sub_wire1(2, 18)    <= sub_wire19(18);
	sub_wire1(2, 19)    <= sub_wire19(19);
	sub_wire1(2, 20)    <= sub_wire19(20);
	sub_wire1(2, 21)    <= sub_wire19(21);
	sub_wire1(2, 22)    <= sub_wire19(22);
	sub_wire1(2, 23)    <= sub_wire19(23);
	sub_wire1(2, 24)    <= sub_wire19(24);
	sub_wire1(2, 25)    <= sub_wire19(25);
	sub_wire1(2, 26)    <= sub_wire19(26);
	sub_wire1(2, 27)    <= sub_wire19(27);
	sub_wire1(2, 28)    <= sub_wire19(28);
	sub_wire1(2, 29)    <= sub_wire19(29);
	sub_wire1(2, 30)    <= sub_wire19(30);
	sub_wire1(2, 31)    <= sub_wire19(31);
	sub_wire1(1, 0)    <= sub_wire20(0);
	sub_wire1(1, 1)    <= sub_wire20(1);
	sub_wire1(1, 2)    <= sub_wire20(2);
	sub_wire1(1, 3)    <= sub_wire20(3);
	sub_wire1(1, 4)    <= sub_wire20(4);
	sub_wire1(1, 5)    <= sub_wire20(5);
	sub_wire1(1, 6)    <= sub_wire20(6);
	sub_wire1(1, 7)    <= sub_wire20(7);
	sub_wire1(1, 8)    <= sub_wire20(8);
	sub_wire1(1, 9)    <= sub_wire20(9);
	sub_wire1(1, 10)    <= sub_wire20(10);
	sub_wire1(1, 11)    <= sub_wire20(11);
	sub_wire1(1, 12)    <= sub_wire20(12);
	sub_wire1(1, 13)    <= sub_wire20(13);
	sub_wire1(1, 14)    <= sub_wire20(14);
	sub_wire1(1, 15)    <= sub_wire20(15);
	sub_wire1(1, 16)    <= sub_wire20(16);
	sub_wire1(1, 17)    <= sub_wire20(17);
	sub_wire1(1, 18)    <= sub_wire20(18);
	sub_wire1(1, 19)    <= sub_wire20(19);
	sub_wire1(1, 20)    <= sub_wire20(20);
	sub_wire1(1, 21)    <= sub_wire20(21);
	sub_wire1(1, 22)    <= sub_wire20(22);
	sub_wire1(1, 23)    <= sub_wire20(23);
	sub_wire1(1, 24)    <= sub_wire20(24);
	sub_wire1(1, 25)    <= sub_wire20(25);
	sub_wire1(1, 26)    <= sub_wire20(26);
	sub_wire1(1, 27)    <= sub_wire20(27);
	sub_wire1(1, 28)    <= sub_wire20(28);
	sub_wire1(1, 29)    <= sub_wire20(29);
	sub_wire1(1, 30)    <= sub_wire20(30);
	sub_wire1(1, 31)    <= sub_wire20(31);
	sub_wire1(0, 0)    <= sub_wire21(0);
	sub_wire1(0, 1)    <= sub_wire21(1);
	sub_wire1(0, 2)    <= sub_wire21(2);
	sub_wire1(0, 3)    <= sub_wire21(3);
	sub_wire1(0, 4)    <= sub_wire21(4);
	sub_wire1(0, 5)    <= sub_wire21(5);
	sub_wire1(0, 6)    <= sub_wire21(6);
	sub_wire1(0, 7)    <= sub_wire21(7);
	sub_wire1(0, 8)    <= sub_wire21(8);
	sub_wire1(0, 9)    <= sub_wire21(9);
	sub_wire1(0, 10)    <= sub_wire21(10);
	sub_wire1(0, 11)    <= sub_wire21(11);
	sub_wire1(0, 12)    <= sub_wire21(12);
	sub_wire1(0, 13)    <= sub_wire21(13);
	sub_wire1(0, 14)    <= sub_wire21(14);
	sub_wire1(0, 15)    <= sub_wire21(15);
	sub_wire1(0, 16)    <= sub_wire21(16);
	sub_wire1(0, 17)    <= sub_wire21(17);
	sub_wire1(0, 18)    <= sub_wire21(18);
	sub_wire1(0, 19)    <= sub_wire21(19);
	sub_wire1(0, 20)    <= sub_wire21(20);
	sub_wire1(0, 21)    <= sub_wire21(21);
	sub_wire1(0, 22)    <= sub_wire21(22);
	sub_wire1(0, 23)    <= sub_wire21(23);
	sub_wire1(0, 24)    <= sub_wire21(24);
	sub_wire1(0, 25)    <= sub_wire21(25);
	sub_wire1(0, 26)    <= sub_wire21(26);
	sub_wire1(0, 27)    <= sub_wire21(27);
	sub_wire1(0, 28)    <= sub_wire21(28);
	sub_wire1(0, 29)    <= sub_wire21(29);
	sub_wire1(0, 30)    <= sub_wire21(30);
	sub_wire1(0, 31)    <= sub_wire21(31);
	result    <= sub_wire22(31 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 21,
		lpm_type => "LPM_MUX",
		lpm_width => 32,
		lpm_widths => 5
	)
	PORT MAP (
		data => sub_wire1,
		sel => sel,
		result => sub_wire22
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "21"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "5"
-- Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL "data0x[31..0]"
-- Retrieval info: USED_PORT: data10x 0 0 32 0 INPUT NODEFVAL "data10x[31..0]"
-- Retrieval info: USED_PORT: data11x 0 0 32 0 INPUT NODEFVAL "data11x[31..0]"
-- Retrieval info: USED_PORT: data12x 0 0 32 0 INPUT NODEFVAL "data12x[31..0]"
-- Retrieval info: USED_PORT: data13x 0 0 32 0 INPUT NODEFVAL "data13x[31..0]"
-- Retrieval info: USED_PORT: data14x 0 0 32 0 INPUT NODEFVAL "data14x[31..0]"
-- Retrieval info: USED_PORT: data15x 0 0 32 0 INPUT NODEFVAL "data15x[31..0]"
-- Retrieval info: USED_PORT: data16x 0 0 32 0 INPUT NODEFVAL "data16x[31..0]"
-- Retrieval info: USED_PORT: data17x 0 0 32 0 INPUT NODEFVAL "data17x[31..0]"
-- Retrieval info: USED_PORT: data18x 0 0 32 0 INPUT NODEFVAL "data18x[31..0]"
-- Retrieval info: USED_PORT: data19x 0 0 32 0 INPUT NODEFVAL "data19x[31..0]"
-- Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL "data1x[31..0]"
-- Retrieval info: USED_PORT: data20x 0 0 32 0 INPUT NODEFVAL "data20x[31..0]"
-- Retrieval info: USED_PORT: data2x 0 0 32 0 INPUT NODEFVAL "data2x[31..0]"
-- Retrieval info: USED_PORT: data3x 0 0 32 0 INPUT NODEFVAL "data3x[31..0]"
-- Retrieval info: USED_PORT: data4x 0 0 32 0 INPUT NODEFVAL "data4x[31..0]"
-- Retrieval info: USED_PORT: data5x 0 0 32 0 INPUT NODEFVAL "data5x[31..0]"
-- Retrieval info: USED_PORT: data6x 0 0 32 0 INPUT NODEFVAL "data6x[31..0]"
-- Retrieval info: USED_PORT: data7x 0 0 32 0 INPUT NODEFVAL "data7x[31..0]"
-- Retrieval info: USED_PORT: data8x 0 0 32 0 INPUT NODEFVAL "data8x[31..0]"
-- Retrieval info: USED_PORT: data9x 0 0 32 0 INPUT NODEFVAL "data9x[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: USED_PORT: sel 0 0 5 0 INPUT NODEFVAL "sel[4..0]"
-- Retrieval info: CONNECT: @data 1 0 32 0 data0x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 10 32 0 data10x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 11 32 0 data11x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 12 32 0 data12x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 13 32 0 data13x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 14 32 0 data14x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 15 32 0 data15x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 16 32 0 data16x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 17 32 0 data17x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 18 32 0 data18x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 19 32 0 data19x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 1 32 0 data1x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 20 32 0 data20x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 2 32 0 data2x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 3 32 0 data3x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 4 32 0 data4x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 5 32 0 data5x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 6 32 0 data6x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 7 32 0 data7x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 8 32 0 data8x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 9 32 0 data9x 0 0 32 0
-- Retrieval info: CONNECT: @sel 0 0 5 0 sel 0 0 5 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ula_mux.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ula_mux.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ula_mux.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ula_mux.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ula_mux_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
